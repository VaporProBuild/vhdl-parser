This is a test VHD file

Remove this file when you use it!!!